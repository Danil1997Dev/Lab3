// dec_test.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module dec_test (
		input  wire  clk_clk,           //        clk.clk
		input  wire  reset_reset_n,     //      reset.reset_n
		input  wire  sem_export_train,  // sem_export.train
		output wire  sem_export_red,    //           .red
		output wire  sem_export_yellow, //           .yellow
		output wire  sem_export_green   //           .green
	);

	wire  [31:0] master_m0_readdata;                        // mm_interconnect_0:master_m0_readdata -> master:avm_readdata
	wire         master_m0_waitrequest;                     // mm_interconnect_0:master_m0_waitrequest -> master:avm_waitrequest
	wire  [31:0] master_m0_address;                         // master:avm_address -> mm_interconnect_0:master_m0_address
	wire         master_m0_read;                            // master:avm_read -> mm_interconnect_0:master_m0_read
	wire   [3:0] master_m0_byteenable;                      // master:avm_byteenable -> mm_interconnect_0:master_m0_byteenable
	wire         master_m0_readdatavalid;                   // mm_interconnect_0:master_m0_readdatavalid -> master:avm_readdatavalid
	wire  [31:0] master_m0_writedata;                       // master:avm_writedata -> mm_interconnect_0:master_m0_writedata
	wire         master_m0_write;                           // master:avm_write -> mm_interconnect_0:master_m0_write
	wire  [31:0] mm_interconnect_0_sem_ctl_slave_readdata;  // sem:ctl_rddata -> mm_interconnect_0:sem_ctl_slave_readdata
	wire   [0:0] mm_interconnect_0_sem_ctl_slave_address;   // mm_interconnect_0:sem_ctl_slave_address -> sem:ctl_addr
	wire         mm_interconnect_0_sem_ctl_slave_read;      // mm_interconnect_0:sem_ctl_slave_read -> sem:ctl_rd
	wire         mm_interconnect_0_sem_ctl_slave_write;     // mm_interconnect_0:sem_ctl_slave_write -> sem:ctl_wr
	wire  [31:0] mm_interconnect_0_sem_ctl_slave_writedata; // mm_interconnect_0:sem_ctl_slave_writedata -> sem:ctl_wrdata
	wire   [1:0] mm_interconnect_0_sem_ram_slave_address;   // mm_interconnect_0:sem_ram_slave_address -> sem:ram_addr
	wire         mm_interconnect_0_sem_ram_slave_write;     // mm_interconnect_0:sem_ram_slave_write -> sem:ram_wr
	wire  [31:0] mm_interconnect_0_sem_ram_slave_writedata; // mm_interconnect_0:sem_ram_slave_writedata -> sem:ram_wrdata
	wire         rst_controller_reset_out_reset;            // rst_controller:reset_out -> [master:reset, mm_interconnect_0:master_clk_reset_reset_bridge_in_reset_reset, sem:clrn]

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (32),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) master (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.avm_address            (master_m0_address),              //        m0.address
		.avm_readdata           (master_m0_readdata),             //          .readdata
		.avm_writedata          (master_m0_writedata),            //          .writedata
		.avm_waitrequest        (master_m0_waitrequest),          //          .waitrequest
		.avm_write              (master_m0_write),                //          .write
		.avm_read               (master_m0_read),                 //          .read
		.avm_byteenable         (master_m0_byteenable),           //          .byteenable
		.avm_readdatavalid      (master_m0_readdatavalid),        //          .readdatavalid
		.avm_burstcount         (),                               // (terminated)
		.avm_begintransfer      (),                               // (terminated)
		.avm_beginbursttransfer (),                               // (terminated)
		.avm_arbiterlock        (),                               // (terminated)
		.avm_lock               (),                               // (terminated)
		.avm_debugaccess        (),                               // (terminated)
		.avm_transactionid      (),                               // (terminated)
		.avm_readid             (8'b00000000),                    // (terminated)
		.avm_writeid            (8'b00000000),                    // (terminated)
		.avm_clken              (),                               // (terminated)
		.avm_response           (2'b00),                          // (terminated)
		.avm_writeresponsevalid (1'b0),                           // (terminated)
		.avm_readresponse       (8'b00000000),                    // (terminated)
		.avm_writeresponse      (8'b00000000)                     // (terminated)
	);

	dec #(
		.m (8)
	) sem (
		.clk        (clk_clk),                                   //      clock.clk
		.clrn       (~rst_controller_reset_out_reset),           // reset_sink.reset_n
		.ctl_rd     (mm_interconnect_0_sem_ctl_slave_read),      //  ctl_slave.read
		.ctl_addr   (mm_interconnect_0_sem_ctl_slave_address),   //           .address
		.ctl_wrdata (mm_interconnect_0_sem_ctl_slave_writedata), //           .writedata
		.ctl_rddata (mm_interconnect_0_sem_ctl_slave_readdata),  //           .readdata
		.ctl_wr     (mm_interconnect_0_sem_ctl_slave_write),     //           .write
		.ram_wr     (mm_interconnect_0_sem_ram_slave_write),     //  ram_slave.write
		.ram_addr   (mm_interconnect_0_sem_ram_slave_address),   //           .address
		.ram_wrdata (mm_interconnect_0_sem_ram_slave_writedata), //           .writedata
		.train      (sem_export_train),                          //        sem.train
		.red        (sem_export_red),                            //           .red
		.yellow     (sem_export_yellow),                         //           .yellow
		.green      (sem_export_green)                           //           .green
	);

	dec_test_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                (clk_clk),                                   //                              clk_0_clk.clk
		.master_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),            // master_clk_reset_reset_bridge_in_reset.reset
		.master_m0_address                            (master_m0_address),                         //                              master_m0.address
		.master_m0_waitrequest                        (master_m0_waitrequest),                     //                                       .waitrequest
		.master_m0_byteenable                         (master_m0_byteenable),                      //                                       .byteenable
		.master_m0_read                               (master_m0_read),                            //                                       .read
		.master_m0_readdata                           (master_m0_readdata),                        //                                       .readdata
		.master_m0_readdatavalid                      (master_m0_readdatavalid),                   //                                       .readdatavalid
		.master_m0_write                              (master_m0_write),                           //                                       .write
		.master_m0_writedata                          (master_m0_writedata),                       //                                       .writedata
		.sem_ctl_slave_address                        (mm_interconnect_0_sem_ctl_slave_address),   //                          sem_ctl_slave.address
		.sem_ctl_slave_write                          (mm_interconnect_0_sem_ctl_slave_write),     //                                       .write
		.sem_ctl_slave_read                           (mm_interconnect_0_sem_ctl_slave_read),      //                                       .read
		.sem_ctl_slave_readdata                       (mm_interconnect_0_sem_ctl_slave_readdata),  //                                       .readdata
		.sem_ctl_slave_writedata                      (mm_interconnect_0_sem_ctl_slave_writedata), //                                       .writedata
		.sem_ram_slave_address                        (mm_interconnect_0_sem_ram_slave_address),   //                          sem_ram_slave.address
		.sem_ram_slave_write                          (mm_interconnect_0_sem_ram_slave_write),     //                                       .write
		.sem_ram_slave_writedata                      (mm_interconnect_0_sem_ram_slave_writedata)  //                                       .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
